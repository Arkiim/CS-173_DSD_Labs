architecture rtl of light_manager_normal is
begin

end architecture rtl;
