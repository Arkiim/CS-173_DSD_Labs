architecture rtl of cycle_manager is
begin

end architecture rtl;
