architecture rtl of light_manager_rush is
begin

end architecture rtl;