architecture rtl of light_manager is
begin

end architecture rtl;
