architecture rtl of bcd_to_7seg is
begin

end architecture rtl;
